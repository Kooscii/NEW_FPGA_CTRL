module i2c_slave(
	//I2C 2-wire
	SDA,
	SCL,
	
	//the data to be analyse
	data,
	command,
	
	//the flag to call recieve successing
	rcv_succ
);

inout SDA;
input SCL;
output [7:0] command;
output[15:0] data;
output rcv_succ;

//I2C slave address
parameter I2C_ADR = 7'h27;

wire SDA_shadow;
wire start_or_stop;
assign SDA_shadow = (~SCL | start_or_stop) ? SDA : SDA_shadow;
assign start_or_stop = ~SCL ? 1'b0 : (SDA ^ SDA_shadow);

reg incycle;
always @(negedge SCL or posedge start_or_stop)
if(start_or_stop)
	incycle <= 1'b0;
	else if(~SDA)
		incycle <= 1'b1;

reg [3:0] bitcnt;  // counts the I2C bits from 7 downto 0, plus an ACK bit
wire bit_DATA = ~bitcnt[3];  // the DATA bits are the first 8 bits sent
wire bit_ACK = bitcnt[3];  // the ACK bit is the 9th bit sent
reg data_phase;

reg[2:0] order;

always @(negedge SCL or negedge incycle)
if(~incycle)	begin
    bitcnt <= 4'h7;  // the bit 7 is received first
    data_phase <= 0;
	 order <= 3'd0;
	end
else	begin
	if(bit_ACK)	begin
		bitcnt <= 4'h7;
		data_phase <= 1;
		order <= order + 1'b1;	//count to 3
		end
		else
			bitcnt <= bitcnt - 4'h1;
	end

wire adr_phase = ~data_phase;
reg adr_match, op_read, got_ACK;
// sample SDA on posedge since the I2C spec specifies as low as 0µs hold-time on negedge
reg SDAr;

always @(posedge SCL)
	SDAr <= SDA;

reg [7:0] mem_1, mem_2, mem_3, mem_4, mem_5,  mem_6;
wire op_write = ~op_read;

always @(negedge SCL or negedge incycle)
if(~incycle)	begin
	got_ACK <= 0;
	adr_match <= 1;
	op_read <= 0;
	end
	else	begin
		if(adr_phase & bitcnt==7 & SDAr!=I2C_ADR[6]) adr_match<=0;
		if(adr_phase & bitcnt==6 & SDAr!=I2C_ADR[5]) adr_match<=0;
		if(adr_phase & bitcnt==5 & SDAr!=I2C_ADR[4]) adr_match<=0;
		if(adr_phase & bitcnt==4 & SDAr!=I2C_ADR[3]) adr_match<=0;
		if(adr_phase & bitcnt==3 & SDAr!=I2C_ADR[2]) adr_match<=0;
		if(adr_phase & bitcnt==2 & SDAr!=I2C_ADR[1]) adr_match<=0;
		if(adr_phase & bitcnt==1 & SDAr!=I2C_ADR[0]) adr_match<=0;
		if(adr_phase & bitcnt==0) op_read <= SDAr;	// 0 slave recieve
		//monitor the ACK to be able to free the bus when the master doesn't ACK during a read operation
		if(bit_ACK) got_ACK <= ~SDAr;	//the BUS released to be pull down
		if((adr_match & bit_DATA & data_phase & op_write) && (order==3'd1)) mem_1[bitcnt] <= SDAr;  // memory write
		if((adr_match & bit_DATA & data_phase & op_write) && (order==3'd2)) mem_2[bitcnt] <= SDAr;  // memory write
		if((adr_match & bit_DATA & data_phase & op_write) && (order==3'd3)) mem_3[bitcnt] <= SDAr;  // memory write
	end
	
//wire mem_bit_low = ~mem_1[bitcnt[2:0]];
//wire SDA_assert_low = adr_match & bit_DATA & data_phase & op_read & mem_bit_low & got_ACK;	//response0
wire SDA_assert_low = adr_match & bit_DATA & data_phase & op_read & got_ACK;	//response0
wire SDA_assert_ACK = adr_match & bit_ACK & (adr_phase | op_write);	//response 1
wire SDA_low = SDA_assert_low | SDA_assert_ACK;
assign SDA = SDA_low ? 1'b0 : 1'bz;

assign command = mem_1; 
assign data = {mem_2,mem_3};

assign rcv_succ = bit_ACK & (order==3'd3) & data_phase;

endmodule